`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/12/02 21:00:21
// Design Name: 
// Module Name: sound_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sound_rom(
	input wire clk,
    input wire [5:0] addr,
    output reg [15:0] data
    );

	 reg [10:0] addr_reg; 

   // body
   always @(posedge clk) 
      addr_reg <= addr;
      
   always @*
      case (addr_reg)
        
         6'h00: data = 16'b0000000100000010; // 
         6'h01: data = 16'b0000001100000100; // 
         6'h02: data = 16'b0000011100001000; // 
         6'h03: data = 16'b0000111100010000; // 
         6'h04: data = 16'b1101111100000000; // 
         6'h05: data = 16'b1101111100000000; // 
         6'h06: data = 16'b1101111100000000; // 
         6'h07: data = 16'b1101111100011110; // 
         6'h08: data = 16'b1101111100000000; // 
         6'h09: data = 16'b1101111100000000; // 
         6'h0a: data = 16'b1101111100000000; // 
         6'h0b: data = 16'b1101111100000000; // 
         6'h0c: data = 16'b0000111100010000; // 
         6'h0d: data = 16'b0000011100001000; // 
         6'h0e: data = 16'b0000001100000100; // 
         6'h0f: data = 16'b0000000100000010; // 
      
         6'h10: data = 16'b0000000100000000; // 
         6'h11: data = 16'b0000001100000000; // 
         6'h12: data = 16'b0000011101000010; // 
         6'h13: data = 16'b0000111101000010; // 
         6'h14: data = 16'b1101111101100110; // 
         6'h15: data = 16'b1101111100100100; // 
         6'h16: data = 16'b1101111100100100; // 
         6'h17: data = 16'b1101111100011000; // 
         6'h18: data = 16'b1101111100011000; // 
         6'h19: data = 16'b1101111100100100; // 
         6'h1a: data = 16'b1101111100100100; // 
         6'h1b: data = 16'b1101111101100110; // 
         6'h1c: data = 16'b0000111101000010; // 
         6'h1d: data = 16'b0000011101000010; // 
         6'h1e: data = 16'b0000001100000000; // 
         6'h1f: data = 16'b0000000100000000; // 

         6'h20: data = 16'b0000000000000000; // 
         6'h21: data = 16'b0000000000000000; // 
         6'h22: data = 16'b0000000000000000; // 
         6'h23: data = 16'b0000000000000000; // 
         6'h24: data = 16'b0000000000000000; // 
         6'h25: data = 16'b0000000000000000; // 
         6'h26: data = 16'b0000000000000000; // 
         6'h27: data = 16'b0000000000000000; // 
         6'h28: data = 16'b0000000000000000; // 
         6'h29: data = 16'b0000000000000000; // 
         6'h2a: data = 16'b0000000000000000; // 
         6'h2b: data = 16'b0000000000000000; // 
         6'h2c: data = 16'b0000000000000000; // 
         6'h2d: data = 16'b0000000000000000; // 
         6'h2e: data = 16'b0000000000000000; // 
         6'h2f: data = 16'b0000000000000000; // 
         
	   endcase

endmodule
