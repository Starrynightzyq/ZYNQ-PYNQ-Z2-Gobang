`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/11/13 19:43:00
// Design Name: 
// Module Name: cursor_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cursor_rom(
	input wire clk,
    input wire [10:0] addr,
    output reg [15:0] data
    );

	 reg [10:0] addr_reg; 

   // body
   always @(posedge clk) 
      addr_reg <= addr;

   always @*
      case (addr_reg)
         //code x00
         11'h000: data = 16'h07E0; // 
         11'h001: data = 16'h1C38; // 
         11'h002: data = 16'h2004; // 
         11'h003: data = 16'h6006; // 
         11'h004: data = 16'h4002; // 
         11'h005: data = 16'hCC33; // 
         11'h006: data = 16'h8C31; // 
         11'h007: data = 16'h8001; // 
         11'h008: data = 16'h8001; // 
         11'h009: data = 16'h8811; // 
         11'h00a: data = 16'hC423; // 
         11'h00b: data = 16'h43C2; // 
         11'h00c: data = 16'h6006; // 
         11'h00d: data = 16'h2004; // 
         11'h00e: data = 16'h1C38; // 
         11'h00f: data = 16'h07E0; // 
         //code x01
         11'h010: data = 16'h07E0; // 
         11'h011: data = 16'h1FF8; // 
         11'h012: data = 16'h3FFC; // 
         11'h013: data = 16'h7FFE; // 
         11'h014: data = 16'h7FFE; // 
         11'h015: data = 16'hF3CF; // 
         11'h016: data = 16'hF3CF; // 
         11'h017: data = 16'hFFFF; // 
         11'h018: data = 16'hFFFF; // 
         11'h019: data = 16'hF7EF; // 
         11'h01a: data = 16'hFBDF; // 
         11'h01b: data = 16'h7C3E; // 
         11'h01c: data = 16'h7FFE; // 
         11'h01d: data = 16'h3FFC; // 
         11'h01e: data = 16'h1FF8; // 
         11'h01f: data = 16'h07E0; // 
         //code x02
         11'h020: data = 16'b1000000000000000; // 
         11'h021: data = 16'b1100000000000000; // 
         11'h022: data = 16'b1010000000000000; // 
         11'h023: data = 16'b1001000000000000; // 
         11'h024: data = 16'b1000100000000000; // 
         11'h025: data = 16'b1000010000000000; // 
         11'h026: data = 16'b1000001000000000; // 
         11'h027: data = 16'b1000000100000000; // 
         11'h028: data = 16'b1000000010000000; // 
         11'h029: data = 16'b1000001111000000; // 
         11'h02a: data = 16'b1001001000000000; // 
         11'h02b: data = 16'b1010100100000000; // 
         11'h02c: data = 16'b1100100100000000; // 
         11'h02d: data = 16'b1000010010000000; // 
         11'h02e: data = 16'b0000010010000000; // 
         11'h02f: data = 16'b0000001100000000; // 
         //code x03
         11'h030: data = 16'b1000000000000000; // 
         11'h031: data = 16'b1100000000000000; // 
         11'h032: data = 16'b1110000000000000; // 
         11'h033: data = 16'b1111000000000000; // 
         11'h034: data = 16'b1111100000000000; // 
         11'h035: data = 16'b1111110000000000; // 
         11'h036: data = 16'b1111111000000000; // 
         11'h037: data = 16'b1111111100000000; // 
         11'h038: data = 16'b1111111110000000; // 
         11'h039: data = 16'b1111111111000000; // 
         11'h03a: data = 16'b1111111000000000; // 
         11'h03b: data = 16'b1110111100000000; // 
         11'h03c: data = 16'b1100111100000000; // 
         11'h03d: data = 16'b1000011110000000; // 
         11'h03e: data = 16'b0000011110000000; // 
         11'h03f: data = 16'b0000001100000000; // 
         //code x04
         11'h040: data = 16'b0000000000000000; // 
         11'h041: data = 16'b0001111111110000; // 
         11'h042: data = 16'b0010000000001000; // 
         11'h043: data = 16'b0010100000101000; // 
         11'h044: data = 16'b0010000000001000; // 
         11'h045: data = 16'b0010000000001000; // 
         11'h046: data = 16'b0010100000101000; // 
         11'h047: data = 16'b0010011111001000; // 
         11'h048: data = 16'b0010000000001000; // 
         11'h049: data = 16'b0001111111110000; // 
         11'h04a: data = 16'b0100000000000100; // 
         11'h04b: data = 16'b0010000000001000; // 
         11'h04c: data = 16'b0011000000011000; // 
         11'h04d: data = 16'b0011000000011000; // 
         11'h04e: data = 16'b0011000000011000; // 
         11'h04f: data = 16'b0000000000000000; // 
         //code x05
         11'h050: data = 16'b0000000000000000; // 
         11'h051: data = 16'b0001111111110000; // 
         11'h052: data = 16'b0011111111111000; // 
         11'h053: data = 16'b0011011111011000; // 
         11'h054: data = 16'b0011111111111000; // 
         11'h055: data = 16'b0011111111111000; // 
         11'h056: data = 16'b0011011111011000; // 
         11'h057: data = 16'b0011100000111000; // 
         11'h058: data = 16'b0011111111111000; // 
         11'h059: data = 16'b0001111111110000; // 
         11'h05a: data = 16'b0100000000000100; // 
         11'h05b: data = 16'b0010000000001000; // 
         11'h05c: data = 16'b0011000000011000; // 
         11'h05d: data = 16'b0011000000011000; // 
         11'h05e: data = 16'b0011000000011000; // 
         11'h05f: data = 16'b0000000000000000; // 
    endcase
endmodule
